module SD_uart_rx #(
    parameter UART_BPS = 'd921600,     //?????????
    parameter CLK_FREQ = 'd20_000_000  //??????
) (
    input wire sys_clk,    //?????50MHz
    input wire sys_rst_n,  //??????
    input wire rx,         //???????????

    output reg [7:0] po_data,  //????????8bit????
    output reg       po_flag   //??????????????????????
);

  //********************************************************************//
  //****************** Parameter and Internal Signal *******************//
  //********************************************************************//
  //localparam    define
  localparam BAUD_CNT_MAX = CLK_FREQ / UART_BPS + 1;
  //reg   define
  reg        rx_reg1;
  reg        rx_reg2;
  reg        rx_reg3;
  reg        start_nedge;
  reg        work_en;
  reg [12:0] baud_cnt;
  reg        bit_flag;
  reg [ 3:0] bit_cnt;
  reg [ 7:0] rx_data;
  reg        rx_flag;
  //********************************************************************//
  //***************************** Main Code ****************************//
  //********************************************************************//
  //???????????????????????????????????????
  //rx_reg1:????????????????????????????1
  always @(posedge sys_clk or negedge sys_rst_n)
    if (sys_rst_n == 1'b0) rx_reg1 <= 1'b1;
    else rx_reg1 <= rx;

  //rx_reg2:????????????????????????????1
  always @(posedge sys_clk or negedge sys_rst_n)
    if (sys_rst_n == 1'b0) rx_reg2 <= 1'b1;
    else rx_reg2 <= rx_reg1;

  //rx_reg3:????????????????????????????????????
  always @(posedge sys_clk or negedge sys_rst_n)
    if (sys_rst_n == 1'b0) rx_reg3 <= 1'b1;
    else rx_reg3 <= rx_reg2;

  //start_nedge:?????????start_nedge??????????????
  always @(posedge sys_clk or negedge sys_rst_n)
    if (sys_rst_n == 1'b0) start_nedge <= 1'b0;
    else if ((~rx_reg2) && (rx_reg3)) start_nedge <= 1'b1;
    else start_nedge <= 1'b0;

  //work_en:?????????????????
  always @(posedge sys_clk or negedge sys_rst_n)
    if (sys_rst_n == 1'b0) work_en <= 1'b0;
    else if (start_nedge == 1'b1) work_en <= 1'b1;
    else if ((bit_cnt == 4'd8) && (bit_flag == 1'b1)) work_en <= 1'b0;

  //baud_cnt:???????????????????0??????BAUD_CNT_MAX - 1
  always @(posedge sys_clk or negedge sys_rst_n)
    if (sys_rst_n == 1'b0) baud_cnt <= 13'b0;
    else if ((baud_cnt == BAUD_CNT_MAX - 1) || (work_en == 1'b0)) baud_cnt <= 13'b0;
    else if (work_en == 1'b1) baud_cnt <= baud_cnt + 1'b1;

  //bit_flag:??baud_cnt????????????????????????????????????
  //?????????????????????????????
  always @(posedge sys_clk or negedge sys_rst_n)
    if (sys_rst_n == 1'b0) bit_flag <= 1'b0;
    else if (baud_cnt == BAUD_CNT_MAX / 2 - 1) bit_flag <= 1'b1;
    else bit_flag <= 1'b0;

  //bit_cnt:?????????????????????8????????????????????????????
  //???????????????????
  always @(posedge sys_clk or negedge sys_rst_n)
    if (sys_rst_n == 1'b0) bit_cnt <= 4'b0;
    else if ((bit_cnt == 4'd8) && (bit_flag == 1'b1)) bit_cnt <= 4'b0;
    else if (bit_flag == 1'b1) bit_cnt <= bit_cnt + 1'b1;

  //rx_data:???????????????
  always @(posedge sys_clk or negedge sys_rst_n)
    if (sys_rst_n == 1'b0) rx_data <= 8'b0;
    else if ((bit_cnt >= 4'd1) && (bit_cnt <= 4'd8) && (bit_flag == 1'b1))
      rx_data <= {rx_reg3, rx_data[7:1]};

  //rx_flag:????????????????rx_flag??????????????
  always @(posedge sys_clk or negedge sys_rst_n)
    if (sys_rst_n == 1'b0) rx_flag <= 1'b0;
    else if ((bit_cnt == 4'd8) && (bit_flag == 1'b1)) rx_flag <= 1'b1;
    else rx_flag <= 1'b0;

  //po_data:?????????8??????????
  always @(posedge sys_clk or negedge sys_rst_n)
    if (sys_rst_n == 1'b0) po_data <= 8'b0;
    else if (rx_flag == 1'b1) po_data <= rx_data;

  //po_flag:??????????????????rx_flag??????????????????po_data?????
  always @(posedge sys_clk or negedge sys_rst_n)
    if (sys_rst_n == 1'b0) po_flag <= 1'b0;
    else po_flag <= rx_flag;

endmodule



////////////////////////////////////////////////////////////////////////
// Author        : EmbedFire
// ?????: ???FPGA???????????????
// ???    : http://www.embedfire.com
// ???    : http://www.firebbs.cn
// ???    : https://fire-stm32.taobao.com
////////////////////////////////////////////////////////////////////////

module Write_sd_init (
    input wire sys_clk,    //?????????,???50MHz
    input wire sys_rst_n,  //?????????,??????????????
    input wire miso,       //?????????????

    output reg cs_n,     //?????????????????
    output reg mosi,     //??????????????
    output reg init_end  //??????????????????
);

  //********************************************************************//
  //****************** Parameter and Internal Signal *******************//
  //********************************************************************//
  //parameter define
  parameter CMD0 = {
    8'h40, 8'h00, 8'h00, 8'h00, 8'h00, 8'h95
  },  //???????
  CMD8 = {
    8'h48, 8'h00, 8'h00, 8'h01, 8'haa, 8'h87
  },  //?????????
  CMD55 = {
    8'h77, 8'h00, 8'h00, 8'h00, 8'h00, 8'hff
  },  //???????????
  ACMD41 = {
    8'h69, 8'h40, 8'h00, 8'h00, 8'h00, 8'hff
  };  //??????
  parameter CNT_WAIT_MAX = 8'd100;  //?????????????????????????
  parameter IDLE = 4'b0000,  //???????
  SEND_CMD0 = 4'b0001,  //CMD0??????????????
  CMD0_ACK = 4'b0011,  //CMD0???????
  SEND_CMD8 = 4'b0010,  //CMD8??????????????
  CMD8_ACK = 4'b0110,  //CMD8???????
  SEND_CMD55 = 4'b0111,  //CMD55??????????????
  CMD55_ACK = 4'b0101,  //CMD55???????
  SEND_ACMD41 = 4'b0100,  //ACMD41??????????????
  ACMD41_ACK = 4'b1100,  //ACMD41???????
  INIT_END = 4'b1101;  //?????????????????

  //reg   define
  reg [ 7:0] cnt_wait;  //????????????????????
  reg [ 3:0] state;  //??????????
  reg [ 7:0] cnt_cmd_bit;  //?????????????????
  reg        miso_dly;  //???????????????????????
  reg        ack_en;  //?????????
  reg [39:0] ack_data;  //???????
  reg [ 7:0] cnt_ack_bit;  //?????????????

  //********************************************************************//
  //***************************** Main Code ****************************//
  //********************************************************************//
  //cnt_wait:????????????????????
  always @(posedge sys_clk or negedge sys_rst_n)
    if (sys_rst_n == 1'b0) cnt_wait <= 8'd0;
    else if (cnt_wait >= CNT_WAIT_MAX) cnt_wait <= CNT_WAIT_MAX;
    else cnt_wait <= cnt_wait + 1'b1;

  //state:???????????????????
  always @(posedge sys_clk or negedge sys_rst_n)
    if (sys_rst_n == 1'b0) state <= IDLE;
    else
      case (state)
        IDLE:
        if (cnt_wait == CNT_WAIT_MAX) state <= SEND_CMD0;
        else state <= state;
        SEND_CMD0:
        if (cnt_cmd_bit == 8'd48) state <= CMD0_ACK;
        else state <= state;
        CMD0_ACK:
        if (cnt_ack_bit == 8'd48)
          if (ack_data[39:32] == 8'h01) state <= SEND_CMD8;
          else state <= SEND_CMD0;
        else state <= state;
        SEND_CMD8:
        if (cnt_cmd_bit == 8'd48) state <= CMD8_ACK;
        else state <= state;
        CMD8_ACK:
        if (cnt_ack_bit == 8'd48)
          if (ack_data[11:8] == 4'b0001) state <= SEND_CMD55;
          else state <= SEND_CMD8;
        else state <= state;
        SEND_CMD55:
        if (cnt_cmd_bit == 8'd48) state <= CMD55_ACK;
        else state <= state;
        CMD55_ACK:
        if (cnt_ack_bit == 8'd48)
          if (ack_data[39:32] == 8'h01) state <= SEND_ACMD41;
          else state <= SEND_CMD55;
        else state <= state;
        SEND_ACMD41:
        if (cnt_cmd_bit == 8'd48) state <= ACMD41_ACK;
        else state <= state;
        ACMD41_ACK:
        if (cnt_ack_bit == 8'd48)
          if (ack_data[39:32] == 8'h00) state <= INIT_END;
          else state <= SEND_CMD55;
        else state <= state;
        INIT_END: state <= state;
        default: state <= IDLE;
      endcase

  //cs_n,mosi,init_end,cnt_cmd_bit
  //?????????????,??????????????,??????????????????,????????????????
  always @(posedge sys_clk or negedge sys_rst_n)
    if (sys_rst_n == 1'b0) begin
      cs_n        <= 1'b1;
      mosi        <= 1'b1;
      init_end    <= 1'b0;
      cnt_cmd_bit <= 8'd0;
    end else
      case (state)
        IDLE: begin
          cs_n        <= 1'b1;
          mosi        <= 1'b1;
          init_end    <= 1'b0;
          cnt_cmd_bit <= 8'd0;
        end
        SEND_CMD0:
        if (cnt_cmd_bit == 8'd48) cnt_cmd_bit <= 8'd0;
        else begin
          cs_n        <= 1'b0;
          mosi        <= CMD0[8'd47-cnt_cmd_bit];
          init_end    <= 1'b0;
          cnt_cmd_bit <= cnt_cmd_bit + 8'd1;
        end
        CMD0_ACK:   if (cnt_ack_bit == 8'd47) cs_n <= 1'b1;
 else cs_n <= 1'b0;
        SEND_CMD8:
        if (cnt_cmd_bit == 8'd48) cnt_cmd_bit <= 8'd0;
        else begin
          cs_n        <= 1'b0;
          mosi        <= CMD8[8'd47-cnt_cmd_bit];
          init_end    <= 1'b0;
          cnt_cmd_bit <= cnt_cmd_bit + 8'd1;
        end
        CMD8_ACK:   if (cnt_ack_bit == 8'd47) cs_n <= 1'b1;
 else cs_n <= 1'b0;
        SEND_CMD55:
        if (cnt_cmd_bit == 8'd48) cnt_cmd_bit <= 8'd0;
        else begin
          cs_n        <= 1'b0;
          mosi        <= CMD55[8'd47-cnt_cmd_bit];
          init_end    <= 1'b0;
          cnt_cmd_bit <= cnt_cmd_bit + 8'd1;
        end
        CMD55_ACK:  if (cnt_ack_bit == 8'd47) cs_n <= 1'b1;
 else cs_n <= 1'b0;
        SEND_ACMD41:
        if (cnt_cmd_bit == 8'd48) cnt_cmd_bit <= 8'd0;
        else begin
          cs_n        <= 1'b0;
          mosi        <= ACMD41[8'd47-cnt_cmd_bit];
          init_end    <= 1'b0;
          cnt_cmd_bit <= cnt_cmd_bit + 8'd1;
        end
        ACMD41_ACK: if (cnt_ack_bit < 8'd47) cs_n <= 1'b0;
 else cs_n <= 1'b1;
        INIT_END: begin
          cs_n     <= 1'b1;
          mosi     <= 1'b1;
          init_end <= 1'b1;
        end
        default: begin
          cs_n <= 1'b1;
          mosi <= 1'b1;
        end
      endcase

  //miso_dly:??????????????????????
  always @(negedge sys_clk or negedge sys_rst_n)
    if (sys_rst_n == 1'b0) miso_dly <= 1'b0;
    else miso_dly <= miso;

  //ack_en:?????????
  always @(negedge sys_clk or negedge sys_rst_n)
    if (sys_rst_n == 1'b0) ack_en <= 1'b0;
    else if (cnt_ack_bit == 8'd47) ack_en <= 1'b0;
    else if ((miso == 1'b0) && (miso_dly == 1'b1) && (cnt_ack_bit == 8'd0)) ack_en <= 1'b1;
    else ack_en <= ack_en;

  //ack_data:???????
  //cnt_ack_bit:?????????????
  always @(negedge sys_clk or negedge sys_rst_n)
    if (sys_rst_n == 1'b0) begin
      ack_data    <=  8'b0;
      cnt_ack_bit <=  8'd0;
    end else if (ack_en == 1'b1) begin
      cnt_ack_bit <= cnt_ack_bit + 8'd1;
      if (cnt_ack_bit < 8'd40) ack_data <= {ack_data[38:0], miso_dly};
      else ack_data <= ack_data;
    end else cnt_ack_bit <= 8'd0;

endmodule

module Write_sd_write (
    input wire        sys_clk,    //?????????,???50MHz
    input wire        sys_rst_n,  //?????????,?????????????
    input wire        miso,       //?????????????
    input wire        wr_en,      //??????????????????
    input wire [31:0] wr_addr,    //???????????????????
    input wire [15:0] wr_data,    //???????????

    output reg  cs_n,     //????????????????
    output reg  mosi,     //??????????????
    output wire wr_busy,  //??????????
    output wire wr_req    //???????????????????
);

  //********************************************************************//
  //****************** Parameter and Internal Signal *******************//
  //********************************************************************//
  //parameter define
  parameter IDLE = 3'b000,  //???????
  SEND_CMD24 = 3'b001,  //??????CMD24?????????????
  CMD24_ACK = 3'b011,  //CMD24???????
  WR_DATA = 3'b010,  //??????????????
  WR_BUSY = 3'b110,  //SD?????????????
  WR_END = 3'b111;  //??????????????
  parameter DATA_NUM = 12'd256;  //???????????????
  parameter BYTE_HEAD = 16'hfffe;  //??????????

  //wire  define
  wire [47:0] cmd_wr;  //??????????????

  //reg   define
  reg  [ 2:0] state;  //??????????
  reg  [ 7:0] cnt_cmd_bit;  //????????????????
  reg         ack_en;  //?????????
  reg  [ 7:0] ack_data;  //???????
  reg  [ 7:0] cnt_ack_bit;  //?????????????
  reg  [11:0] cnt_data_num;  //???????????????
  reg  [ 3:0] cnt_data_bit;  //??????????????
  reg  [ 7:0] busy_data;  //????????????
  reg  [ 2:0] cnt_end;  //???????????????????
  reg         miso_dly;  //??????????????????????

  //********************************************************************//
  //***************************** Main Code ****************************//
  //********************************************************************//
  //wr_busy:??????????
  assign wr_busy = (state != IDLE) ? 1'b1 : 1'b0;

  //wr_req:???????????????????
  assign wr_req  = ((cnt_data_num <= DATA_NUM - 1'b1) && (cnt_data_bit == 4'd15)) ? 1'b1 : 1'b0;

  //cmd_wr:??????????????
  assign cmd_wr  = {8'h58, wr_addr, 8'hff};

  //miso_dly:??????????????????????
  always @(negedge sys_clk or negedge sys_rst_n)
    if (sys_rst_n == 1'b0) miso_dly <= 1'b0;
    else miso_dly <= miso;

  //ack_en:?????????
  always @(negedge sys_clk or negedge sys_rst_n)
    if (sys_rst_n == 1'b0) ack_en <= 1'b0;
    else if (cnt_ack_bit == 8'd15) ack_en <= 1'b0;
    else if ((state == CMD24_ACK) && (miso == 1'b0) && (miso_dly == 1'b1) && (cnt_ack_bit == 8'd0))
      ack_en <= 1'b1;
    else ack_en <= ack_en;

  //ack_data:???????
  //cnt_ack_bit:?????????????
  always @(negedge sys_clk or negedge sys_rst_n)
    if (sys_rst_n == 1'b0) begin
      ack_data    <=  8'b0;
      cnt_ack_bit <=  8'd0;
    end else if (ack_en == 1'b1) begin
      cnt_ack_bit <= cnt_ack_bit + 8'd1;
      if (cnt_ack_bit < 8'd8) ack_data <= {ack_data[6:0], miso_dly};
      else ack_data <= ack_data;
    end else cnt_ack_bit <= 8'd0;

  //busy_data:????????????
  always @(negedge sys_clk or negedge sys_rst_n)
    if (sys_rst_n == 1'b0) busy_data <= 8'd0;
    else if (state == WR_BUSY) busy_data <= {busy_data[6:0], miso};
    else busy_data <= 8'd0;

  //state:???????????????????
  always @(posedge sys_clk or negedge sys_rst_n)
    if (sys_rst_n == 1'b0) state <= IDLE;
    else
      case (state)
        IDLE:
        if (wr_en == 1'b1) state <= SEND_CMD24;
        else state <= state;
        SEND_CMD24:
        if (cnt_cmd_bit == 8'd47) state <= CMD24_ACK;
        else state <= state;
        CMD24_ACK:
        if (cnt_ack_bit == 8'd15)
          if (ack_data == 8'h00) state <= WR_DATA;
          else state <= SEND_CMD24;
        else state <= state;
        WR_DATA:
        if ((cnt_data_num == (DATA_NUM + 1'b1)) && (cnt_data_bit == 4'd15)) state <= WR_BUSY;
        else state <= state;
        WR_BUSY:
        if (busy_data == 8'hff) state <= WR_END;
        else state <= state;
        WR_END:
        if (cnt_end == 3'd7) state <= IDLE;
        else state <= state;
        default: state <= IDLE;
      endcase

  //cs_n:????????????????
  always @(posedge sys_clk or negedge sys_rst_n)
    if (sys_rst_n == 1'b0) cs_n <= 1'b1;
    else if (cnt_end == 3'd7) cs_n <= 1'b1;
    else if (wr_en == 1'b1) cs_n <= 1'b0;
    else cs_n <= cs_n;

  //cnt_cmd_bit:????????????????
  always @(posedge sys_clk or negedge sys_rst_n)
    if (sys_rst_n == 1'b0) cnt_cmd_bit <= 8'd0;
    else if (state == SEND_CMD24) cnt_cmd_bit <= cnt_cmd_bit + 8'd1;
    else cnt_cmd_bit <= 8'd0;

  //mosi:??????????????
  always @(posedge sys_clk or negedge sys_rst_n)
    if (sys_rst_n == 1'b0) mosi <= 1'b1;
    else if (state == SEND_CMD24) mosi <= cmd_wr[8'd47-cnt_cmd_bit];
    else if (state == WR_DATA)
      if (cnt_data_num == 12'd0) mosi <= BYTE_HEAD[15-cnt_data_bit];
      else if ((cnt_data_num >= 12'd1) && (cnt_data_num <= DATA_NUM))
        mosi <= wr_data[15-cnt_data_bit];
      else mosi <= 1'b1;
    else mosi <= 1'b1;

  //cnt_data_bit:??????????????
  always @(posedge sys_clk or negedge sys_rst_n)
    if (sys_rst_n == 1'b0) cnt_data_bit <= 4'd0;
    else if (state == WR_DATA) cnt_data_bit <= cnt_data_bit + 4'd1;
    else cnt_data_bit <= 4'd0;

  //cnt_data_num:???????????????
  always @(posedge sys_clk or negedge sys_rst_n)
    if (sys_rst_n == 1'b0) cnt_data_num <= 12'd0;
    else if (state == WR_DATA)
      if (cnt_data_bit == 4'd15) cnt_data_num <= cnt_data_num + 12'd1;
      else cnt_data_num <= cnt_data_num;
    else cnt_data_num <= 12'd0;

  //cnt_end:???????????????????
  always @(posedge sys_clk or negedge sys_rst_n)
    if (sys_rst_n == 1'b0) cnt_end <= 3'd0;
    else if (state == WR_END) cnt_end <= cnt_end + 3'd1;
    else cnt_end <= 3'd0;

endmodule


////////////////////////////////////////////////////////////////////////
// Author        : EmbedFire
// ?????: ???FPGA??????????????
// ???    : http://www.embedfire.com
// ???    : http://www.firebbs.cn
// ???    : https://fire-stm32.taobao.com
////////////////////////////////////////////////////////////////////////

module Write_sd_Control (
    input  wire        sys_clk,     //?????????,???50MHz
    input  wire        sys_rst_n,   //?????????,?????????????
    //SD???????????
    input  wire        sd_miso,     //?????????????
    output wire        sd_clk,      //SD??????????????
    output reg         sd_cs_n,     //?????????????
    output reg         sd_mosi,     //??????????????
    //??SD???????????
    input  wire        wr_en,       //??????????????????
    input  wire [31:0] wr_addr,     //???????????????????
    input  wire [15:0] wr_data,     //???????????
    output wire        wr_busy,     //??????????
    output wire        wr_req,      //???????????????????
    //??SD???????????
    input  wire        rd_en,       //?????????????????
    input  wire [31:0] rd_addr,     //???????????????????
    output wire        rd_busy,     //??????????
    output wire        rd_data_en,  //?????????????????
    output wire [15:0] rd_data,     //???????????

    output wire init_end  //SD?????????????
);

  //********************************************************************//
  //****************** Parameter and Internal Signal *******************//
  //********************************************************************//
  //wire define
  wire init_cs_n;  //???????????????????
  wire init_mosi;  //????????????????????????????
  wire wr_cs_n;  //???????????????????
  wire wr_mosi;  //????????????????????????????
  wire rd_cs_n;  //???????????????????
  wire rd_mosi;  //????????????????????????????

  //********************************************************************//
  //***************************** Main Code ****************************//
  //********************************************************************//
  //sd_clk:SD??????????????
  assign sd_clk = !sys_clk;

  //SD?????????????
  always @(*)
    if (init_end == 1'b0) begin
      sd_cs_n <= init_cs_n;
      sd_mosi <= init_mosi;
    end else if (wr_busy == 1'b1) begin
      sd_cs_n <= wr_cs_n;
      sd_mosi <= wr_mosi;
    end else if (rd_busy == 1'b1) begin
      sd_cs_n <= rd_cs_n;
      sd_mosi <= rd_mosi;
    end else begin
      sd_cs_n <= 1'b1;
      sd_mosi <= 1'b1;
    end

  //********************************************************************//
  //************************** Instantiation ***************************//
  //********************************************************************//
  //------------- sd_init_inst -------------
  Write_sd_init sd_init_inst (
      .sys_clk  (sys_clk),    //?????????,???50MHz
      .sys_rst_n(sys_rst_n),  //?????????,?????????????
      .miso     (sd_miso),    //?????????????

      .cs_n    (init_cs_n),  //????????????????
      .mosi    (init_mosi),  //??????????????
      .init_end(init_end)    //?????????????????
  );

  //------------- sd_write_inst -------------
  Write_sd_write sd_write_inst (
      .sys_clk  (sys_clk),            //?????????,???50MHz
      .sys_rst_n(sys_rst_n),          //?????????,?????????????
      .miso     (sd_miso),            //?????????????
      .wr_en    (wr_en && init_end),  //??????????????????
      .wr_addr  (wr_addr),            //???????????????????
      .wr_data  (wr_data),            //???????????

      .cs_n   (wr_cs_n),  //????????????????
      .mosi   (wr_mosi),  //??????????????
      .wr_busy(wr_busy),  //??????????
      .wr_req (wr_req)    //???????????????????
  );

endmodule


////////////////////////////////////////////////////////////////////////
// Author        : EmbedFire
// ?????: ???FPGA???????????????
// ???    : http://www.embedfire.com
// ???    : http://www.firebbs.cn
// ???    : https://fire-stm32.taobao.com
////////////////////////////////////////////////////////////////////////

module SDDataWriter (
    //??????
    input  wire        sys_clk,    //?????????,???50MHz
    input  wire        sys_rst_n,  //?????????,?????????????
    //??????
    input  wire        rx_flag,    //??fifo?????????????
    input  wire [ 7:0] rx_data,    //??fifo????????
    //SD???????
    input  wire        sd_miso,    //?????????????
    output wire        sd_clk,     //SD??????????????
    output wire        sd_cs_n,    //?????????????
    output wire        sd_mosi,    //??????????????
    //??SD????
    inout  wire        wr_en,      //??????????????????
    input  wire [31:0] wr_addr,    //???????????????????
    inout  wire [15:0] wr_data,    //???????????
    output wire        wr_busy,    //??????????
    output wire        wr_req      //???????????????????
);

  //********************************************************************//
  //****************** Parameter and Internal Signal *******************//
  //********************************************************************//
  //parameter define
  parameter DATA_NUM = 12'd256;  //???????????
  parameter SECTOR_ADDR = 32'd1000;  //???????????????
  parameter CNT_WAIT_MAX = 16'd60000;  //??fifo?????????????????????????????

  //wire  define
  wire [11:0] wr_fifo_data_num;  //??fifo???????????????
  wire        wr_busy_fall;  //sd?????????????????
  wire        rd_busy_fall;  //sd?????????????????
  wire        init_end;  //?????SD???
  //reg   define
  reg         wr_busy_dly;  //sd?????????????????????????????
  reg         rd_busy_dly;  //sd?????????????????????????????
  reg         send_data_en;  //?????????????????????????
  reg  [15:0] cnt_wait;  //??fifo????????????????
  reg  [11:0] send_data_num;  //?????????????????????
  reg         rd_fifo_rd_en;


  wire        rd_data_en;  //sd??????????????????????
  wire [15:0] rd_data;  //sd????????????????
  wire        rd_busy;  //sd???????????????????
  reg         rd_en;  //sd?????????????
  wire [31:0] rd_addr;  //sd???????????????
  reg         tx_flag;  //??fifo?????????????
  wire [ 7:0] tx_data;  //??fifo????????
  //********************************************************************//
  //***************************** Main Code ****************************//
  //********************************************************************//
  //wr_en:sd??????????????
  assign wr_en = (((wr_fifo_data_num == (DATA_NUM)) && (init_end == 1'b1))) ? 1'b1 : 1'b0;

  //wr_busy_dly:sd?????????????????????????????
  always @(posedge sys_clk or negedge sys_rst_n)
    if (sys_rst_n == 1'b0) wr_busy_dly <= 1'b0;
    else wr_busy_dly <= wr_busy;

  //wr_busy_fall:sd?????????????????
  assign wr_busy_fall = ((wr_busy == 1'b0) && (wr_busy_dly == 1'b1)) ? 1'b1 : 1'b0;

  //rd_en:sd?????????????
  always @(posedge sys_clk or negedge sys_rst_n)
    if (sys_rst_n == 1'b0) rd_en <= 1'b0;
    else if (wr_busy_fall == 1'b1) rd_en <= 1'b1;
    else rd_en <= 1'b0;

  //rd_addr:sd???????????????
  assign rd_addr = SECTOR_ADDR;

  //rd_busy_dly:sd?????????????????????????????
  always @(posedge sys_clk or negedge sys_rst_n)
    if (sys_rst_n == 1'b0) rd_busy_dly <= 1'b0;
    else rd_busy_dly <= rd_busy;

  //rd_busy_fall:sd?????????????????
  assign rd_busy_fall = ((rd_busy == 1'b0) && (rd_busy_dly == 1'b1)) ? 1'b1 : 1'b0;

  //send_data_en:?????????????????????????
  always @(posedge sys_clk or negedge sys_rst_n)
    if (sys_rst_n == 1'b0) send_data_en <= 1'b0;
    else if ((send_data_num == (DATA_NUM * 2) - 1'b1) && (cnt_wait == CNT_WAIT_MAX - 1'b1))
      send_data_en <= 1'b0;
    else if (rd_busy_fall == 1'b1) send_data_en <= 1'b1;
    else send_data_en <= send_data_en;

  //cnt_wait:??fifo????????????????
  always @(posedge sys_clk or negedge sys_rst_n)
    if (sys_rst_n == 1'b0) cnt_wait <= 16'd0;
    else if (send_data_en == 1'b1)
      if (cnt_wait == CNT_WAIT_MAX) cnt_wait <= 16'd0;
      else cnt_wait <= cnt_wait + 1'b1;
    else cnt_wait <= 16'd0;

  //send_data_num:?????????????????????
  always @(posedge sys_clk or negedge sys_rst_n)
    if (sys_rst_n == 1'b0) send_data_num <= 12'd0;
    else if (send_data_en == 1'b1)
      if (cnt_wait == CNT_WAIT_MAX) send_data_num <= send_data_num + 1'b1;
      else send_data_num <= send_data_num;
    else send_data_num <= 12'd0;

  //rd_fifo_rd_en:??fifo???????????????
  always @(posedge sys_clk or negedge sys_rst_n)
    if (sys_rst_n == 1'b0) rd_fifo_rd_en <= 1'b0;
    else if (cnt_wait == (CNT_WAIT_MAX - 1'b1)) rd_fifo_rd_en <= 1'b1;
    else rd_fifo_rd_en <= 1'b0;

  //tx_flag:??fifo?????????????
  always @(posedge sys_clk or negedge sys_rst_n)
    if (sys_rst_n == 1'b0) tx_flag <= 1'b0;
    else tx_flag <= rd_fifo_rd_en;

  //********************************************************************//
  //************************** Instantiation ***************************//
  //********************************************************************//
  //------------- fifo_wr_data_inst -------------
  wr_fifo fifo_wr_data_inst (
      .rst   (~sys_rst_n),  //??��
      .wr_clk(sys_clk),     //????��?????????
      .wr_en (rx_flag),     //????��?????????
      .din   (rx_data),     //��??????

      .full         (),
      .empty        (),
      .rd_clk       (sys_clk),          //??????????????
      .rd_en        (wr_req),           //??????????????
      .dout         (wr_data),          //????????
      .rd_data_count(wr_fifo_data_num)  //fifo??????????????????
  );
  ila_0 FIFODebug (
      .clk   (sys_clk),
      .probe0(~sys_rst_n),
      .probe1(sys_clk),     //SD卡时钟信�????
      .probe2(rx_flag),     //片�?�信�????
      .probe3(wr_req)
  );
  Write_sd_Control SDControl (
      .sys_clk  (sys_clk),   //?????????,???50MHz
      .sys_rst_n(sys_rst_n), //?????????,???????????????

      .sd_miso(sd_miso),  //?????????????
      .sd_clk (sd_clk),   //SD????????????????
      .sd_cs_n(sd_cs_n),  //???????????????
      .sd_mosi(sd_mosi),  //??????????????

      .wr_en  (wr_en),    //????????????????????
      .wr_addr(wr_addr),  //?????????????????????
      .wr_data(wr_data),  //?????????????
      .wr_busy(wr_busy),  //??????????
      .wr_req (wr_req),   //?????????????????????

      .init_end(init_end)  //SD??????
  );

endmodule

module WriteAddressChange (

    input  wire        AddOnce,
    input  wire        sys_rst_n,           //?????????,?????????????
    input  wire [31:0] StartWriterAddress,  //sd???????????????
    output reg  [31:0] NowWriterAddress     //sd???????????????

);
  //assign  NowWriterAddress = 
  always @(posedge AddOnce or negedge sys_rst_n) begin
    if (!sys_rst_n) begin
      NowWriterAddress <= StartWriterAddress;
    end else begin
      NowWriterAddress <= NowWriterAddress + 32'b1;
    end
  end

endmodule

module WriteSDCardByUART (
    //input  wire Button,
    input  wire sys_clk,    //?????????,???50MHz
    input  wire sys_rst_n,  //?????????,?????????????
    input  wire rx,         //?????????????????
    //    input   wire            SaveToNext  ,   //????????????????????????????????????????????????????
    input  wire sd_miso,    //?????????????
    output wire sd_clk,     //SD??????????????
    output wire sd_cs_n,    //?????????????
    output wire sd_mosi,    //??????????????
    output wire tx

);

  //********************************************************************//
  //****************** Parameter and Internal Signal *******************//
  //********************************************************************//
  //parameter define
  parameter SaveDataAddress = 32'h100;  //??fifo?????????????????????????????

  //wire  define
  wire        rx_flag;  //??fifo?????????????
  wire [ 7:0] rx_data;  //??fifo????????
  wire        wr_req;  //sd????????????
  wire        wr_busy;  //sd??????????????????
  wire        wr_en;  //sd??????????????
  wire [15:0] wr_data;  //sd????????
  wire        rd_data_en;  //sd?????????????????????
  wire [15:0] rd_data;  //sd???????????????
  wire        rd_busy;  //sd??????????????????
  wire        rd_en;  //sd?????????????
  wire [31:0] rd_addr;  //sd???????????????
  wire        tx_flag;  //??fifo?????????????
  wire [ 7:0] tx_data;  //??fifo????????
  wire        locked;  //??????????
  wire        init_end;  //SD?????????????
  wire        CLK_OUT2;
  wire [31:0] WriterAddress;

  //rst_n:???????,???????????


  //------------- SD_uart_rx_inst -------------
  SD_uart_rx SD_uart_rx_inst (
      .sys_clk  (sys_clk),    //?????50Mhz
      .sys_rst_n(sys_rst_n),  //??????
      .rx       (rx),         //???????????

      .po_data(rx_data),  //?????????????????
      .po_flag(rx_flag)   //????????????????????????????
  );
  uart_tx uart_tx_inst (
      .sys_clk  (sys_clk),    //input             sys_clk
      .sys_rst_n(sys_rst_n),  //input             sys_rst_n
      .pi_data  (rx_data),    //input     [7:0]   pi_data
      .pi_flag  (rx_flag),    //input             pi_flag

      .tx(tx)  //output            tx
  );

  WriteAddressChange getTheRealAddress (
      .AddOnce           (wr_en),
      .sys_rst_n         (sys_rst_n),        //?????????,?????????????
      .StartWriterAddress(SaveDataAddress),
      .NowWriterAddress  (WriterAddress)

  );
  SDDataWriter SDControl (
      .sys_clk  (sys_clk),   //?????????,???50MHz
      .sys_rst_n(sys_rst_n), //?????????,?????????????

      .rx_flag(rx_flag),  //??fifo?????????????
      .rx_data(rx_data),  //??fifo????????

      .sd_miso(sd_miso),  //?????????????
      .sd_clk (sd_clk),   //SD??????????????
      .sd_cs_n(sd_cs_n),  //?????????????
      .sd_mosi(sd_mosi),  //??????????????

      .wr_en  (wr_en),          //??????????????????
      .wr_addr(WriterAddress),  //???????????????????
      .wr_data(wr_data),        //???????????
      .wr_busy(wr_busy),        //??????????
      .wr_req (wr_req)          //???????????????????
  );
endmodule
