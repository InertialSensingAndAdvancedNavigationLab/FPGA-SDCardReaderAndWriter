module WriteAddressChange (
    input  wire        AddOnce,
    input  wire        sys_rst_n,           //?????????,?????????????
    output reg  [31:0] NowWriterAddress     //sd???????????????
);

  parameter SaveDataAddress = 32'h0;  //??fifo?????????????????????????????
  //assign  NowWriterAddress = 
  always @(posedge AddOnce or negedge sys_rst_n) begin
    if (!sys_rst_n) begin
      NowWriterAddress <= SaveDataAddress;
    end else begin
      NowWriterAddress <= NowWriterAddress + 32'b1;
    end
  end

endmodule

module WriteSDCardByUART (
    input  wire sys_clk,    //?????????,???50MHz
    input  wire sys_rst,  //?????????,?????????????
    input  wire rx,         //?????????????????
    //    input   wire            SaveToNext  ,   //????????????????????????????????????????????????????
    input  wire sd_miso,    //?????????????
    output wire sd_clk,     //SD??????????????
    output wire sd_cs_n,    //?????????????
    output wire sd_mosi,    //??????????????
    // Debug
    output wire tx

);

  //********************************************************************//
  //****************** Parameter and Internal Signal *******************//
  //********************************************************************//
  //parameter define

  //wire  define
  wire        rx_flag;  //??fifo?????????????
  wire [ 7:0] rx_data;  //??fifo????????
  wire        wr_req;  //sd????????????
  wire        wr_busy;  //sd??????????????????
  wire        wr_en;  //sd??????????????
  wire [15:0] wr_data;  //sd????????
  wire        rd_data_en;  //sd?????????????????????
  wire [15:0] rd_data;  //sd???????????????
  wire        rd_busy;  //sd??????????????????
  wire        rd_en;  //sd?????????????
  wire [31:0] rd_addr;  //sd???????????????
  wire        tx_flag;  //??fifo?????????????
  wire [ 7:0] tx_data;  //??fifo????????
  wire [31:0] WriterAddress;
  // 将rst信号取反得到rst_n信号
  wire sys_rst_n;
  assign sys_rst_n=~sys_rst;
  //------------- SDUartRX_inst -------------
  SDUartRX SDUartInput (
      .sys_clk  (sys_clk),    //?????50Mhz
      .sys_rst_n(sys_rst_n),  //??????
      .rx       (rx),         //???????????

      .po_data(rx_data),  //?????????????????
      .po_flag(rx_flag)   //????????????????????????????
  );
  // Debug Uart Output
  SDUartTX DebugTxOutput (
      .sys_clk  (sys_clk),    //input             sys_clk
      .sys_rst_n(sys_rst_n),  //input             sys_rst_n
      .pi_data  (wr_data),    //input     [7:0]   pi_data
      .pi_flag  (wr_en),    //input             pi_flag

      .tx(tx)  //output            tx
  );

  WriteAddressChange getTheRealAddress (
      .AddOnce           (wr_en),
      .sys_rst_n         (sys_rst_n),
      .NowWriterAddress  (WriterAddress)

  );
  SDDataInput SDControl (
      .sys_clk  (sys_clk),   //?????????,???50MHz
      .sys_rst_n(sys_rst_n), //?????????,?????????????

      .rx_flag(rx_flag),  //??fifo?????????????
      .rx_data(rx_data),  //??fifo????????

      .sd_miso(sd_miso),  //?????????????
      .sd_clk (sd_clk),   //SD??????????????
      .sd_cs_n(sd_cs_n),  //?????????????
      .sd_mosi(sd_mosi),  //??????????????

      .wr_en  (wr_en),          //??????????????????
      .wr_addr(WriterAddress),  //???????????????????
      .wr_data(wr_data),        //???????????
      .wr_busy(wr_busy),        //??????????
      .wr_req (wr_req)          //???????????????????
  );
endmodule
